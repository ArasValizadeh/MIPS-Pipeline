module ShiftLeft2(
    output [31:0] result,
    input [31:0] input1
);
assign result = input1 << 2;
endmodule
